magic
tech scmos
timestamp 1332627727
<< end >>
