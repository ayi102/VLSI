magic
tech scmos
timestamp 1332529218
<< polysilicon >>
rect -9 20 -7 22
rect -9 18 -2 20
rect -43 16 -41 18
rect -28 16 -26 18
rect -4 16 -2 18
rect 11 19 13 22
rect 11 17 33 19
rect 11 16 13 17
rect 31 16 33 17
rect 46 16 48 18
rect -43 -8 -41 12
rect -28 -8 -26 12
rect -4 -8 -2 12
rect 11 -8 13 12
rect 31 -8 33 12
rect 46 -8 48 12
rect -43 -16 -41 -12
rect -28 -14 -26 -12
rect -4 -16 -2 -12
rect 11 -14 13 -12
rect 31 -14 33 -12
rect 46 -14 48 -12
rect -43 -18 -2 -16
<< ndiffusion >>
rect -45 -12 -43 -8
rect -41 -12 -28 -8
rect -26 -12 -25 -8
rect -6 -12 -4 -8
rect -2 -12 11 -8
rect 13 -12 14 -8
rect 29 -12 31 -8
rect 33 -12 46 -8
rect 48 -12 49 -8
<< pdiffusion >>
rect -45 12 -43 16
rect -41 12 -37 16
rect -33 12 -28 16
rect -26 12 -25 16
rect -6 12 -4 16
rect -2 12 2 16
rect 6 12 11 16
rect 13 12 14 16
rect 29 12 31 16
rect 33 12 37 16
rect 41 12 46 16
rect 48 12 49 16
<< metal1 >>
rect -48 69 -37 74
rect -48 54 -44 69
rect -98 50 -44 54
rect -98 -16 -94 50
rect 2 16 6 20
rect 37 16 41 20
rect -49 8 -45 12
rect -25 8 -21 12
rect -10 8 -6 12
rect 14 8 18 12
rect 25 8 29 12
rect 49 8 53 12
rect -49 4 -21 8
rect -10 4 18 8
rect 25 4 53 8
rect -49 -8 -45 4
rect -37 -4 -33 0
rect -22 -4 -18 0
rect -10 -8 -6 4
rect 2 -4 6 0
rect 17 -4 21 0
rect 25 -8 29 4
rect 37 -4 41 0
rect 52 -4 56 0
rect -65 -16 -61 -10
rect 14 -16 18 -12
rect 49 -16 53 -12
rect -98 -20 53 -16
<< metal2 >>
rect -44 112 60 116
rect -44 101 -40 112
rect -57 23 25 27
rect -57 15 -10 19
rect -14 8 -10 15
rect 21 8 25 23
rect 56 0 60 112
rect -14 -4 -10 0
rect -14 -8 60 -4
<< ntransistor >>
rect -43 -12 -41 -8
rect -28 -12 -26 -8
rect -4 -12 -2 -8
rect 11 -12 13 -8
rect 31 -12 33 -8
rect 46 -12 48 -8
<< ptransistor >>
rect -43 12 -41 16
rect -28 12 -26 16
rect -4 12 -2 16
rect 11 12 13 16
rect 31 12 33 16
rect 46 12 48 16
<< polycontact >>
rect -41 -4 -37 0
rect -26 -4 -22 0
rect -2 -4 2 0
rect 13 -4 17 0
rect 33 -4 37 0
rect 48 -4 52 0
<< ndcontact >>
rect -49 -12 -45 -8
rect -25 -12 -21 -8
rect -10 -12 -6 -8
rect 14 -12 18 -8
rect 25 -12 29 -8
rect 49 -12 53 -8
<< pdcontact >>
rect -49 12 -45 16
rect -37 12 -33 16
rect -25 12 -21 16
rect -10 12 -6 16
rect 2 12 6 16
rect 14 12 18 16
rect 25 12 29 16
rect 37 12 41 16
rect 49 12 53 16
<< m2contact >>
rect -44 97 -40 101
rect -14 4 -10 8
rect 21 4 25 8
rect -18 -4 -14 0
rect 56 -4 60 0
use 3-bitNAND 3-bitNAND_0
timestamp 1332529218
transform 1 0 -144 0 1 23
box 54 -33 107 13
<< end >>
