magic
tech scmos
timestamp 1333126486
<< polysilicon >>
rect -33 -28 -8 -26
rect -33 -40 -31 -28
rect -18 -32 -16 -30
rect -10 -32 -8 -28
rect -2 -28 23 -26
rect -2 -32 0 -28
rect 6 -32 8 -30
rect -33 -54 -31 -44
rect -18 -46 -16 -36
rect -22 -48 -16 -46
rect -22 -52 -20 -48
rect -22 -54 -16 -52
rect -33 -82 -31 -58
rect -18 -66 -16 -54
rect -10 -66 -8 -36
rect -2 -66 0 -36
rect 6 -46 8 -36
rect 21 -40 23 -28
rect 47 -28 72 -26
rect 47 -40 49 -28
rect 62 -32 64 -30
rect 70 -32 72 -28
rect 78 -28 103 -26
rect 78 -32 80 -28
rect 86 -32 88 -30
rect 6 -48 12 -46
rect 10 -52 12 -48
rect 6 -54 12 -52
rect 6 -66 8 -54
rect 21 -55 23 -44
rect 47 -54 49 -44
rect 62 -46 64 -36
rect 58 -48 64 -46
rect 58 -52 60 -48
rect 58 -54 64 -52
rect 21 -61 23 -59
rect 47 -60 49 -58
rect 62 -66 64 -54
rect 70 -66 72 -36
rect 78 -66 80 -36
rect 86 -46 88 -36
rect 101 -40 103 -28
rect 86 -48 92 -46
rect 90 -52 92 -48
rect 86 -54 92 -52
rect 86 -66 88 -54
rect 101 -55 103 -44
rect 101 -61 103 -59
rect -18 -72 -16 -70
rect -10 -72 -8 -70
rect -2 -74 0 -70
rect 6 -72 8 -70
rect 62 -72 64 -70
rect 70 -72 72 -70
rect -25 -76 25 -74
rect 78 -76 80 -70
rect 86 -72 88 -70
rect -25 -82 -23 -76
rect -5 -82 -3 -80
rect 3 -82 5 -80
rect 23 -82 25 -76
rect 31 -78 80 -76
rect 31 -82 33 -78
rect 47 -82 49 -80
rect 58 -82 60 -80
rect 73 -82 75 -80
rect -33 -98 -31 -86
rect -25 -98 -23 -86
rect -5 -98 -3 -86
rect 3 -98 5 -86
rect 23 -98 25 -86
rect 31 -98 33 -86
rect -33 -106 -31 -102
rect -25 -104 -23 -102
rect -5 -106 -3 -102
rect -33 -108 -3 -106
rect 3 -106 5 -102
rect 23 -104 25 -102
rect 31 -106 33 -102
rect 3 -108 33 -106
rect 47 -108 49 -86
rect 58 -108 60 -86
rect 73 -108 75 -86
rect 47 -114 49 -112
rect 58 -114 60 -112
rect 73 -114 75 -112
<< ndiffusion >>
rect -34 -58 -33 -54
rect -31 -58 -30 -54
rect 20 -59 21 -55
rect 23 -59 24 -55
rect 46 -58 47 -54
rect 49 -58 50 -54
rect 100 -59 101 -55
rect 103 -59 104 -55
rect -19 -70 -18 -66
rect -16 -70 -15 -66
rect -11 -70 -10 -66
rect -8 -70 -2 -66
rect 0 -70 1 -66
rect 5 -70 6 -66
rect 8 -70 9 -66
rect 61 -70 62 -66
rect 64 -70 65 -66
rect 69 -70 70 -66
rect 72 -70 78 -66
rect 80 -70 81 -66
rect 85 -70 86 -66
rect 88 -70 89 -66
rect -34 -86 -33 -82
rect -31 -86 -25 -82
rect -23 -86 -22 -82
rect -6 -86 -5 -82
rect -3 -86 3 -82
rect 5 -86 6 -82
rect 22 -86 23 -82
rect 25 -86 31 -82
rect 33 -86 34 -82
rect 46 -86 47 -82
rect 49 -86 58 -82
rect 60 -86 73 -82
rect 75 -86 76 -82
<< pdiffusion >>
rect -19 -36 -18 -32
rect -16 -36 -15 -32
rect -11 -36 -10 -32
rect -8 -36 -7 -32
rect -3 -36 -2 -32
rect 0 -36 1 -32
rect 5 -36 6 -32
rect 8 -36 9 -32
rect -34 -44 -33 -40
rect -31 -44 -30 -40
rect 61 -36 62 -32
rect 64 -36 65 -32
rect 69 -36 70 -32
rect 72 -36 73 -32
rect 77 -36 78 -32
rect 80 -36 81 -32
rect 85 -36 86 -32
rect 88 -36 89 -32
rect 20 -44 21 -40
rect 23 -44 24 -40
rect 46 -44 47 -40
rect 49 -44 50 -40
rect 100 -44 101 -40
rect 103 -44 104 -40
rect -34 -102 -33 -98
rect -31 -102 -30 -98
rect -26 -102 -25 -98
rect -23 -102 -22 -98
rect -6 -102 -5 -98
rect -3 -102 -2 -98
rect 2 -102 3 -98
rect 5 -102 6 -98
rect 22 -102 23 -98
rect 25 -102 26 -98
rect 30 -102 31 -98
rect 33 -102 34 -98
rect 46 -112 47 -108
rect 49 -112 53 -108
rect 57 -112 58 -108
rect 60 -112 61 -108
rect 65 -112 73 -108
rect 75 -112 76 -108
<< metal1 >>
rect -48 -28 108 -24
rect -48 -106 -44 -28
rect -38 -40 -34 -28
rect -7 -32 -3 -28
rect -23 -40 -19 -36
rect -15 -40 -11 -36
rect 1 -40 5 -36
rect -15 -44 5 -40
rect 9 -40 13 -36
rect 24 -40 28 -28
rect 42 -40 46 -28
rect 73 -32 77 -28
rect 57 -40 61 -36
rect 65 -40 69 -36
rect 81 -40 85 -36
rect 65 -44 85 -40
rect 89 -40 93 -36
rect 104 -40 108 -28
rect -41 -51 -37 -47
rect -30 -54 -26 -44
rect -7 -54 -3 -52
rect -15 -58 -3 -54
rect 16 -55 20 -44
rect 27 -52 31 -48
rect 39 -51 43 -47
rect 50 -54 54 -44
rect 73 -54 77 -52
rect -38 -74 -34 -58
rect -23 -66 -19 -62
rect -15 -66 -11 -58
rect 9 -66 13 -62
rect 1 -74 5 -70
rect 24 -74 28 -59
rect 65 -58 77 -54
rect 96 -55 100 -44
rect 107 -52 111 -48
rect 42 -74 46 -58
rect 57 -66 61 -62
rect 65 -66 69 -58
rect 89 -66 93 -62
rect 81 -74 85 -70
rect 104 -74 108 -59
rect -38 -78 108 -74
rect -38 -82 -34 -78
rect -10 -82 -6 -78
rect 18 -82 22 -78
rect 42 -82 46 -78
rect -22 -90 -18 -86
rect 6 -90 10 -86
rect 34 -90 38 -86
rect -38 -94 -18 -90
rect -10 -94 10 -90
rect 18 -91 38 -90
rect 18 -94 43 -91
rect -38 -98 -34 -94
rect -22 -98 -18 -94
rect -10 -98 -6 -94
rect 6 -98 10 -94
rect 18 -98 22 -94
rect 34 -95 43 -94
rect 50 -93 54 -88
rect 65 -92 69 -87
rect 34 -98 38 -95
rect 76 -100 80 -86
rect -30 -106 -26 -102
rect -2 -106 2 -102
rect 26 -106 30 -102
rect 53 -104 80 -100
rect -48 -110 37 -106
rect 53 -108 57 -104
rect 76 -108 80 -104
rect 33 -116 37 -110
rect 42 -116 46 -112
rect 61 -116 65 -112
rect 33 -120 78 -116
<< metal2 >>
rect -23 -48 -19 -44
rect 9 -48 13 -44
rect 31 -48 35 -47
rect -23 -52 -7 -48
rect -3 -51 35 -48
rect 57 -48 61 -44
rect 89 -48 93 -44
rect -3 -52 31 -51
rect 57 -52 73 -48
rect 77 -52 93 -48
rect -19 -62 9 -58
rect 61 -62 89 -58
rect -18 -106 -14 -94
rect 10 -99 14 -94
rect 50 -99 54 -97
rect 10 -102 54 -99
rect 65 -106 69 -96
rect -18 -111 69 -106
<< ntransistor >>
rect -33 -58 -31 -54
rect 21 -59 23 -55
rect 47 -58 49 -54
rect 101 -59 103 -55
rect -18 -70 -16 -66
rect -10 -70 -8 -66
rect -2 -70 0 -66
rect 6 -70 8 -66
rect 62 -70 64 -66
rect 70 -70 72 -66
rect 78 -70 80 -66
rect 86 -70 88 -66
rect -33 -86 -31 -82
rect -25 -86 -23 -82
rect -5 -86 -3 -82
rect 3 -86 5 -82
rect 23 -86 25 -82
rect 31 -86 33 -82
rect 47 -86 49 -82
rect 58 -86 60 -82
rect 73 -86 75 -82
<< ptransistor >>
rect -18 -36 -16 -32
rect -10 -36 -8 -32
rect -2 -36 0 -32
rect 6 -36 8 -32
rect -33 -44 -31 -40
rect 62 -36 64 -32
rect 70 -36 72 -32
rect 78 -36 80 -32
rect 86 -36 88 -32
rect 21 -44 23 -40
rect 47 -44 49 -40
rect 101 -44 103 -40
rect -33 -102 -31 -98
rect -25 -102 -23 -98
rect -5 -102 -3 -98
rect 3 -102 5 -98
rect 23 -102 25 -98
rect 31 -102 33 -98
rect 47 -112 49 -108
rect 58 -112 60 -108
rect 73 -112 75 -108
<< polycontact >>
rect -37 -51 -33 -47
rect -26 -51 -22 -47
rect 12 -52 16 -48
rect 23 -52 27 -48
rect 43 -51 47 -47
rect 54 -51 58 -47
rect 92 -52 96 -48
rect 103 -52 107 -48
rect 43 -95 47 -91
rect 54 -92 58 -88
rect 69 -91 73 -87
<< ndcontact >>
rect -38 -58 -34 -54
rect -30 -58 -26 -54
rect 16 -59 20 -55
rect 24 -59 28 -55
rect 42 -58 46 -54
rect 50 -58 54 -54
rect 96 -59 100 -55
rect 104 -59 108 -55
rect -23 -70 -19 -66
rect -15 -70 -11 -66
rect 1 -70 5 -66
rect 9 -70 13 -66
rect 57 -70 61 -66
rect 65 -70 69 -66
rect 81 -70 85 -66
rect 89 -70 93 -66
rect -38 -86 -34 -82
rect -22 -86 -18 -82
rect -10 -86 -6 -82
rect 6 -86 10 -82
rect 18 -86 22 -82
rect 34 -86 38 -82
rect 42 -86 46 -82
rect 76 -86 80 -82
<< pdcontact >>
rect -23 -36 -19 -32
rect -15 -36 -11 -32
rect -7 -36 -3 -32
rect 1 -36 5 -32
rect 9 -36 13 -32
rect -38 -44 -34 -40
rect -30 -44 -26 -40
rect 57 -36 61 -32
rect 65 -36 69 -32
rect 73 -36 77 -32
rect 81 -36 85 -32
rect 89 -36 93 -32
rect 16 -44 20 -40
rect 24 -44 28 -40
rect 42 -44 46 -40
rect 50 -44 54 -40
rect 96 -44 100 -40
rect 104 -44 108 -40
rect -38 -102 -34 -98
rect -30 -102 -26 -98
rect -22 -102 -18 -98
rect -10 -102 -6 -98
rect -2 -102 2 -98
rect 6 -102 10 -98
rect 18 -102 22 -98
rect 26 -102 30 -98
rect 34 -102 38 -98
rect 42 -112 46 -108
rect 53 -112 57 -108
rect 61 -112 65 -108
rect 76 -112 80 -108
<< m2contact >>
rect -23 -44 -19 -40
rect 9 -44 13 -40
rect 57 -44 61 -40
rect 89 -44 93 -40
rect -7 -52 -3 -48
rect 35 -51 39 -47
rect 73 -52 77 -48
rect -23 -62 -19 -58
rect 9 -62 13 -58
rect 57 -62 61 -58
rect 89 -62 93 -58
rect -18 -94 -14 -90
rect 10 -94 14 -90
rect 50 -97 54 -93
rect 65 -96 69 -92
use 2-bitXOR 2-bitXOR_0
timestamp 1332627727
transform 1 0 14 0 1 23
box 0 0 1 1
use 2-bitXOR 2-bitXOR_1
timestamp 1332627727
transform 1 0 -27 0 1 -55
box 0 0 1 1
use 2-bitXOR 2-bitXOR_2
timestamp 1332627727
transform 1 0 53 0 1 -55
box 0 0 1 1
<< labels >>
rlabel metal1 3 -76 3 -76 1 GND
rlabel metal1 -5 -27 -5 -27 5 VDD
rlabel metal1 75 -56 75 -56 1 SUM
rlabel metal1 109 -50 109 -50 7 CIN
rlabel metal1 29 -50 29 -50 1 B
rlabel metal1 -39 -49 -39 -49 3 A
rlabel metal1 78 -99 78 -99 1 COUT
<< end >>
