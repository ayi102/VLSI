magic
tech scmos
timestamp 1333733533
<< polysilicon >>
rect -33 -28 -8 -26
rect -33 -40 -31 -28
rect -18 -32 -16 -30
rect -10 -32 -8 -28
rect -2 -28 23 -26
rect -2 -32 0 -28
rect 6 -32 8 -30
rect -33 -54 -31 -44
rect -18 -46 -16 -36
rect -22 -48 -16 -46
rect -22 -52 -20 -48
rect -22 -54 -16 -52
rect -33 -82 -31 -58
rect -18 -66 -16 -54
rect -10 -66 -8 -36
rect -2 -66 0 -36
rect 6 -46 8 -36
rect 21 -40 23 -28
rect 47 -28 72 -26
rect 47 -40 49 -28
rect 62 -32 64 -30
rect 70 -32 72 -28
rect 78 -28 103 -26
rect 78 -32 80 -28
rect 86 -32 88 -30
rect 6 -48 12 -46
rect 10 -52 12 -48
rect 6 -54 12 -52
rect 6 -66 8 -54
rect 21 -55 23 -44
rect 47 -54 49 -44
rect 62 -46 64 -36
rect 58 -48 64 -46
rect 58 -52 60 -48
rect 58 -54 64 -52
rect 21 -61 23 -59
rect 47 -60 49 -58
rect 62 -66 64 -54
rect 70 -66 72 -36
rect 78 -66 80 -36
rect 86 -46 88 -36
rect 101 -40 103 -28
rect 86 -48 92 -46
rect 90 -52 92 -48
rect 86 -54 92 -52
rect 86 -66 88 -54
rect 101 -55 103 -44
rect 101 -61 103 -59
rect -18 -72 -16 -70
rect -10 -72 -8 -70
rect -2 -74 0 -70
rect 6 -72 8 -70
rect 62 -72 64 -70
rect 70 -72 72 -70
rect -25 -76 25 -74
rect 78 -76 80 -70
rect 86 -72 88 -70
rect -25 -82 -23 -76
rect -5 -82 -3 -80
rect 3 -82 5 -80
rect 23 -82 25 -76
rect 31 -78 80 -76
rect 31 -82 33 -78
rect 47 -82 49 -80
rect 58 -82 60 -80
rect 73 -82 75 -80
rect -33 -98 -31 -86
rect -25 -98 -23 -86
rect -5 -98 -3 -86
rect 3 -98 5 -86
rect 23 -98 25 -86
rect 31 -98 33 -86
rect -33 -106 -31 -102
rect -25 -104 -23 -102
rect -5 -106 -3 -102
rect -33 -108 -3 -106
rect 3 -106 5 -102
rect 23 -104 25 -102
rect 31 -106 33 -102
rect 3 -108 33 -106
rect 47 -108 49 -86
rect 58 -108 60 -86
rect 73 -108 75 -86
rect 47 -114 49 -112
rect 58 -114 60 -112
rect 73 -114 75 -112
rect -33 -119 -8 -117
rect -33 -131 -31 -119
rect -18 -123 -16 -121
rect -10 -123 -8 -119
rect -2 -119 23 -117
rect -2 -123 0 -119
rect 6 -123 8 -121
rect -33 -145 -31 -135
rect -18 -137 -16 -127
rect -22 -139 -16 -137
rect -22 -143 -20 -139
rect -22 -145 -16 -143
rect -33 -173 -31 -149
rect -18 -157 -16 -145
rect -10 -157 -8 -127
rect -2 -157 0 -127
rect 6 -137 8 -127
rect 21 -131 23 -119
rect 47 -119 72 -117
rect 47 -131 49 -119
rect 62 -123 64 -121
rect 70 -123 72 -119
rect 78 -119 103 -117
rect 78 -123 80 -119
rect 86 -123 88 -121
rect 6 -139 12 -137
rect 10 -143 12 -139
rect 6 -145 12 -143
rect 6 -157 8 -145
rect 21 -146 23 -135
rect 47 -145 49 -135
rect 62 -137 64 -127
rect 58 -139 64 -137
rect 58 -143 60 -139
rect 58 -145 64 -143
rect 21 -152 23 -150
rect 47 -151 49 -149
rect 62 -157 64 -145
rect 70 -157 72 -127
rect 78 -157 80 -127
rect 86 -137 88 -127
rect 101 -131 103 -119
rect 86 -139 92 -137
rect 90 -143 92 -139
rect 86 -145 92 -143
rect 86 -157 88 -145
rect 101 -146 103 -135
rect 101 -152 103 -150
rect -18 -163 -16 -161
rect -10 -163 -8 -161
rect -2 -165 0 -161
rect 6 -163 8 -161
rect 62 -163 64 -161
rect 70 -163 72 -161
rect -25 -167 25 -165
rect 78 -167 80 -161
rect 86 -163 88 -161
rect -25 -173 -23 -167
rect -5 -173 -3 -171
rect 3 -173 5 -171
rect 23 -173 25 -167
rect 31 -169 80 -167
rect 31 -173 33 -169
rect 47 -173 49 -171
rect 58 -173 60 -171
rect 73 -173 75 -171
rect -33 -189 -31 -177
rect -25 -189 -23 -177
rect -5 -189 -3 -177
rect 3 -189 5 -177
rect 23 -189 25 -177
rect 31 -189 33 -177
rect -33 -197 -31 -193
rect -25 -195 -23 -193
rect -5 -197 -3 -193
rect -33 -199 -3 -197
rect 3 -197 5 -193
rect 23 -195 25 -193
rect 31 -197 33 -193
rect 3 -199 33 -197
rect 47 -199 49 -177
rect 58 -199 60 -177
rect 73 -199 75 -177
rect 47 -205 49 -203
rect 58 -205 60 -203
rect 73 -205 75 -203
rect -33 -211 -8 -209
rect -33 -223 -31 -211
rect -18 -215 -16 -213
rect -10 -215 -8 -211
rect -2 -211 23 -209
rect -2 -215 0 -211
rect 6 -215 8 -213
rect -33 -237 -31 -227
rect -18 -229 -16 -219
rect -22 -231 -16 -229
rect -22 -235 -20 -231
rect -22 -237 -16 -235
rect -33 -265 -31 -241
rect -18 -249 -16 -237
rect -10 -249 -8 -219
rect -2 -249 0 -219
rect 6 -229 8 -219
rect 21 -223 23 -211
rect 47 -211 72 -209
rect 47 -223 49 -211
rect 62 -215 64 -213
rect 70 -215 72 -211
rect 78 -211 103 -209
rect 78 -215 80 -211
rect 86 -215 88 -213
rect 6 -231 12 -229
rect 10 -235 12 -231
rect 6 -237 12 -235
rect 6 -249 8 -237
rect 21 -238 23 -227
rect 47 -237 49 -227
rect 62 -229 64 -219
rect 58 -231 64 -229
rect 58 -235 60 -231
rect 58 -237 64 -235
rect 21 -244 23 -242
rect 47 -243 49 -241
rect 62 -249 64 -237
rect 70 -249 72 -219
rect 78 -249 80 -219
rect 86 -229 88 -219
rect 101 -223 103 -211
rect 86 -231 92 -229
rect 90 -235 92 -231
rect 86 -237 92 -235
rect 86 -249 88 -237
rect 101 -238 103 -227
rect 101 -244 103 -242
rect -18 -255 -16 -253
rect -10 -255 -8 -253
rect -2 -257 0 -253
rect 6 -255 8 -253
rect 62 -255 64 -253
rect 70 -255 72 -253
rect -25 -259 25 -257
rect 78 -259 80 -253
rect 86 -255 88 -253
rect -25 -265 -23 -259
rect -5 -265 -3 -263
rect 3 -265 5 -263
rect 23 -265 25 -259
rect 31 -261 80 -259
rect 31 -265 33 -261
rect 47 -265 49 -263
rect 58 -265 60 -263
rect 73 -265 75 -263
rect -33 -281 -31 -269
rect -25 -281 -23 -269
rect -5 -281 -3 -269
rect 3 -281 5 -269
rect 23 -281 25 -269
rect 31 -281 33 -269
rect -33 -289 -31 -285
rect -25 -287 -23 -285
rect -5 -289 -3 -285
rect -33 -291 -3 -289
rect 3 -289 5 -285
rect 23 -287 25 -285
rect 31 -289 33 -285
rect 3 -291 33 -289
rect 47 -291 49 -269
rect 58 -291 60 -269
rect 73 -291 75 -269
rect 47 -297 49 -295
rect 58 -297 60 -295
rect 73 -297 75 -295
rect -33 -303 -8 -301
rect -33 -315 -31 -303
rect -18 -307 -16 -305
rect -10 -307 -8 -303
rect -2 -303 23 -301
rect -2 -307 0 -303
rect 6 -307 8 -305
rect -33 -329 -31 -319
rect -18 -321 -16 -311
rect -22 -323 -16 -321
rect -22 -327 -20 -323
rect -22 -329 -16 -327
rect -33 -357 -31 -333
rect -18 -341 -16 -329
rect -10 -341 -8 -311
rect -2 -341 0 -311
rect 6 -321 8 -311
rect 21 -315 23 -303
rect 47 -303 72 -301
rect 47 -315 49 -303
rect 62 -307 64 -305
rect 70 -307 72 -303
rect 78 -303 103 -301
rect 78 -307 80 -303
rect 86 -307 88 -305
rect 6 -323 12 -321
rect 10 -327 12 -323
rect 6 -329 12 -327
rect 6 -341 8 -329
rect 21 -330 23 -319
rect 47 -329 49 -319
rect 62 -321 64 -311
rect 58 -323 64 -321
rect 58 -327 60 -323
rect 58 -329 64 -327
rect 21 -336 23 -334
rect 47 -335 49 -333
rect 62 -341 64 -329
rect 70 -341 72 -311
rect 78 -341 80 -311
rect 86 -321 88 -311
rect 101 -315 103 -303
rect 86 -323 92 -321
rect 90 -327 92 -323
rect 86 -329 92 -327
rect 86 -341 88 -329
rect 101 -330 103 -319
rect 101 -336 103 -334
rect -18 -347 -16 -345
rect -10 -347 -8 -345
rect -2 -349 0 -345
rect 6 -347 8 -345
rect 62 -347 64 -345
rect 70 -347 72 -345
rect -25 -351 25 -349
rect 78 -351 80 -345
rect 86 -347 88 -345
rect -25 -357 -23 -351
rect -5 -357 -3 -355
rect 3 -357 5 -355
rect 23 -357 25 -351
rect 31 -353 80 -351
rect 31 -357 33 -353
rect 47 -357 49 -355
rect 58 -357 60 -355
rect 73 -357 75 -355
rect -33 -373 -31 -361
rect -25 -373 -23 -361
rect -5 -373 -3 -361
rect 3 -373 5 -361
rect 23 -373 25 -361
rect 31 -373 33 -361
rect -33 -381 -31 -377
rect -25 -379 -23 -377
rect -5 -381 -3 -377
rect -33 -383 -3 -381
rect 3 -381 5 -377
rect 23 -379 25 -377
rect 31 -381 33 -377
rect 3 -383 33 -381
rect 47 -383 49 -361
rect 58 -383 60 -361
rect 73 -383 75 -361
rect 47 -389 49 -387
rect 58 -389 60 -387
rect 73 -389 75 -387
<< ndiffusion >>
rect -34 -58 -33 -54
rect -31 -58 -30 -54
rect 20 -59 21 -55
rect 23 -59 24 -55
rect 46 -58 47 -54
rect 49 -58 50 -54
rect 100 -59 101 -55
rect 103 -59 104 -55
rect -19 -70 -18 -66
rect -16 -70 -15 -66
rect -11 -70 -10 -66
rect -8 -70 -2 -66
rect 0 -70 1 -66
rect 5 -70 6 -66
rect 8 -70 9 -66
rect 61 -70 62 -66
rect 64 -70 65 -66
rect 69 -70 70 -66
rect 72 -70 78 -66
rect 80 -70 81 -66
rect 85 -70 86 -66
rect 88 -70 89 -66
rect -34 -86 -33 -82
rect -31 -86 -25 -82
rect -23 -86 -22 -82
rect -6 -86 -5 -82
rect -3 -86 3 -82
rect 5 -86 6 -82
rect 22 -86 23 -82
rect 25 -86 31 -82
rect 33 -86 34 -82
rect 46 -86 47 -82
rect 49 -86 58 -82
rect 60 -86 73 -82
rect 75 -86 76 -82
rect -34 -149 -33 -145
rect -31 -149 -30 -145
rect 20 -150 21 -146
rect 23 -150 24 -146
rect 46 -149 47 -145
rect 49 -149 50 -145
rect 100 -150 101 -146
rect 103 -150 104 -146
rect -19 -161 -18 -157
rect -16 -161 -15 -157
rect -11 -161 -10 -157
rect -8 -161 -2 -157
rect 0 -161 1 -157
rect 5 -161 6 -157
rect 8 -161 9 -157
rect 61 -161 62 -157
rect 64 -161 65 -157
rect 69 -161 70 -157
rect 72 -161 78 -157
rect 80 -161 81 -157
rect 85 -161 86 -157
rect 88 -161 89 -157
rect -34 -177 -33 -173
rect -31 -177 -25 -173
rect -23 -177 -22 -173
rect -6 -177 -5 -173
rect -3 -177 3 -173
rect 5 -177 6 -173
rect 22 -177 23 -173
rect 25 -177 31 -173
rect 33 -177 34 -173
rect 46 -177 47 -173
rect 49 -177 58 -173
rect 60 -177 73 -173
rect 75 -177 76 -173
rect -34 -241 -33 -237
rect -31 -241 -30 -237
rect 20 -242 21 -238
rect 23 -242 24 -238
rect 46 -241 47 -237
rect 49 -241 50 -237
rect 100 -242 101 -238
rect 103 -242 104 -238
rect -19 -253 -18 -249
rect -16 -253 -15 -249
rect -11 -253 -10 -249
rect -8 -253 -2 -249
rect 0 -253 1 -249
rect 5 -253 6 -249
rect 8 -253 9 -249
rect 61 -253 62 -249
rect 64 -253 65 -249
rect 69 -253 70 -249
rect 72 -253 78 -249
rect 80 -253 81 -249
rect 85 -253 86 -249
rect 88 -253 89 -249
rect -34 -269 -33 -265
rect -31 -269 -25 -265
rect -23 -269 -22 -265
rect -6 -269 -5 -265
rect -3 -269 3 -265
rect 5 -269 6 -265
rect 22 -269 23 -265
rect 25 -269 31 -265
rect 33 -269 34 -265
rect 46 -269 47 -265
rect 49 -269 58 -265
rect 60 -269 73 -265
rect 75 -269 76 -265
rect -34 -333 -33 -329
rect -31 -333 -30 -329
rect 20 -334 21 -330
rect 23 -334 24 -330
rect 46 -333 47 -329
rect 49 -333 50 -329
rect 100 -334 101 -330
rect 103 -334 104 -330
rect -19 -345 -18 -341
rect -16 -345 -15 -341
rect -11 -345 -10 -341
rect -8 -345 -2 -341
rect 0 -345 1 -341
rect 5 -345 6 -341
rect 8 -345 9 -341
rect 61 -345 62 -341
rect 64 -345 65 -341
rect 69 -345 70 -341
rect 72 -345 78 -341
rect 80 -345 81 -341
rect 85 -345 86 -341
rect 88 -345 89 -341
rect -34 -361 -33 -357
rect -31 -361 -25 -357
rect -23 -361 -22 -357
rect -6 -361 -5 -357
rect -3 -361 3 -357
rect 5 -361 6 -357
rect 22 -361 23 -357
rect 25 -361 31 -357
rect 33 -361 34 -357
rect 46 -361 47 -357
rect 49 -361 58 -357
rect 60 -361 73 -357
rect 75 -361 76 -357
<< pdiffusion >>
rect -19 -36 -18 -32
rect -16 -36 -15 -32
rect -11 -36 -10 -32
rect -8 -36 -7 -32
rect -3 -36 -2 -32
rect 0 -36 1 -32
rect 5 -36 6 -32
rect 8 -36 9 -32
rect -34 -44 -33 -40
rect -31 -44 -30 -40
rect 61 -36 62 -32
rect 64 -36 65 -32
rect 69 -36 70 -32
rect 72 -36 73 -32
rect 77 -36 78 -32
rect 80 -36 81 -32
rect 85 -36 86 -32
rect 88 -36 89 -32
rect 20 -44 21 -40
rect 23 -44 24 -40
rect 46 -44 47 -40
rect 49 -44 50 -40
rect 100 -44 101 -40
rect 103 -44 104 -40
rect -34 -102 -33 -98
rect -31 -102 -30 -98
rect -26 -102 -25 -98
rect -23 -102 -22 -98
rect -6 -102 -5 -98
rect -3 -102 -2 -98
rect 2 -102 3 -98
rect 5 -102 6 -98
rect 22 -102 23 -98
rect 25 -102 26 -98
rect 30 -102 31 -98
rect 33 -102 34 -98
rect 46 -112 47 -108
rect 49 -112 53 -108
rect 57 -112 58 -108
rect 60 -112 61 -108
rect 65 -112 73 -108
rect 75 -112 76 -108
rect -19 -127 -18 -123
rect -16 -127 -15 -123
rect -11 -127 -10 -123
rect -8 -127 -7 -123
rect -3 -127 -2 -123
rect 0 -127 1 -123
rect 5 -127 6 -123
rect 8 -127 9 -123
rect -34 -135 -33 -131
rect -31 -135 -30 -131
rect 61 -127 62 -123
rect 64 -127 65 -123
rect 69 -127 70 -123
rect 72 -127 73 -123
rect 77 -127 78 -123
rect 80 -127 81 -123
rect 85 -127 86 -123
rect 88 -127 89 -123
rect 20 -135 21 -131
rect 23 -135 24 -131
rect 46 -135 47 -131
rect 49 -135 50 -131
rect 100 -135 101 -131
rect 103 -135 104 -131
rect -34 -193 -33 -189
rect -31 -193 -30 -189
rect -26 -193 -25 -189
rect -23 -193 -22 -189
rect -6 -193 -5 -189
rect -3 -193 -2 -189
rect 2 -193 3 -189
rect 5 -193 6 -189
rect 22 -193 23 -189
rect 25 -193 26 -189
rect 30 -193 31 -189
rect 33 -193 34 -189
rect 46 -203 47 -199
rect 49 -203 53 -199
rect 57 -203 58 -199
rect 60 -203 61 -199
rect 65 -203 73 -199
rect 75 -203 76 -199
rect -19 -219 -18 -215
rect -16 -219 -15 -215
rect -11 -219 -10 -215
rect -8 -219 -7 -215
rect -3 -219 -2 -215
rect 0 -219 1 -215
rect 5 -219 6 -215
rect 8 -219 9 -215
rect -34 -227 -33 -223
rect -31 -227 -30 -223
rect 61 -219 62 -215
rect 64 -219 65 -215
rect 69 -219 70 -215
rect 72 -219 73 -215
rect 77 -219 78 -215
rect 80 -219 81 -215
rect 85 -219 86 -215
rect 88 -219 89 -215
rect 20 -227 21 -223
rect 23 -227 24 -223
rect 46 -227 47 -223
rect 49 -227 50 -223
rect 100 -227 101 -223
rect 103 -227 104 -223
rect -34 -285 -33 -281
rect -31 -285 -30 -281
rect -26 -285 -25 -281
rect -23 -285 -22 -281
rect -6 -285 -5 -281
rect -3 -285 -2 -281
rect 2 -285 3 -281
rect 5 -285 6 -281
rect 22 -285 23 -281
rect 25 -285 26 -281
rect 30 -285 31 -281
rect 33 -285 34 -281
rect 46 -295 47 -291
rect 49 -295 53 -291
rect 57 -295 58 -291
rect 60 -295 61 -291
rect 65 -295 73 -291
rect 75 -295 76 -291
rect -19 -311 -18 -307
rect -16 -311 -15 -307
rect -11 -311 -10 -307
rect -8 -311 -7 -307
rect -3 -311 -2 -307
rect 0 -311 1 -307
rect 5 -311 6 -307
rect 8 -311 9 -307
rect -34 -319 -33 -315
rect -31 -319 -30 -315
rect 61 -311 62 -307
rect 64 -311 65 -307
rect 69 -311 70 -307
rect 72 -311 73 -307
rect 77 -311 78 -307
rect 80 -311 81 -307
rect 85 -311 86 -307
rect 88 -311 89 -307
rect 20 -319 21 -315
rect 23 -319 24 -315
rect 46 -319 47 -315
rect 49 -319 50 -315
rect 100 -319 101 -315
rect 103 -319 104 -315
rect -34 -377 -33 -373
rect -31 -377 -30 -373
rect -26 -377 -25 -373
rect -23 -377 -22 -373
rect -6 -377 -5 -373
rect -3 -377 -2 -373
rect 2 -377 3 -373
rect 5 -377 6 -373
rect 22 -377 23 -373
rect 25 -377 26 -373
rect 30 -377 31 -373
rect 33 -377 34 -373
rect 46 -387 47 -383
rect 49 -387 53 -383
rect 57 -387 58 -383
rect 60 -387 61 -383
rect 65 -387 73 -383
rect 75 -387 76 -383
<< metal1 >>
rect -48 -28 108 -24
rect -48 -106 -44 -28
rect -38 -40 -34 -28
rect -7 -32 -3 -28
rect -23 -40 -19 -36
rect -15 -40 -11 -36
rect 1 -40 5 -36
rect -15 -44 5 -40
rect 9 -40 13 -36
rect 24 -40 28 -28
rect 42 -40 46 -28
rect 73 -32 77 -28
rect 57 -40 61 -36
rect 65 -40 69 -36
rect 81 -40 85 -36
rect 65 -44 85 -40
rect 89 -40 93 -36
rect 104 -40 108 -28
rect -41 -51 -37 -47
rect -30 -54 -26 -44
rect -7 -54 -3 -52
rect -15 -58 -3 -54
rect 16 -55 20 -44
rect 27 -52 31 -48
rect 39 -51 43 -47
rect 50 -54 54 -44
rect 73 -54 77 -52
rect -38 -74 -34 -58
rect -23 -66 -19 -62
rect -15 -66 -11 -58
rect 9 -66 13 -62
rect 1 -74 5 -70
rect 24 -74 28 -59
rect 65 -58 77 -54
rect 96 -55 100 -44
rect 107 -52 111 -48
rect 42 -74 46 -58
rect 57 -66 61 -62
rect 65 -66 69 -58
rect 89 -66 93 -62
rect 81 -74 85 -70
rect 104 -74 108 -59
rect -38 -78 108 -74
rect -38 -82 -34 -78
rect -10 -82 -6 -78
rect 18 -82 22 -78
rect 42 -82 46 -78
rect -22 -90 -18 -86
rect 6 -90 10 -86
rect 34 -90 38 -86
rect -38 -94 -18 -90
rect -10 -94 10 -90
rect 18 -91 38 -90
rect 18 -94 43 -91
rect -38 -98 -34 -94
rect -22 -98 -18 -94
rect -10 -98 -6 -94
rect 6 -98 10 -94
rect 18 -98 22 -94
rect 34 -95 43 -94
rect 50 -93 54 -88
rect 65 -92 69 -87
rect 76 -90 80 -86
rect 34 -98 38 -95
rect 76 -94 115 -90
rect 76 -100 80 -94
rect -30 -106 -26 -102
rect -2 -106 2 -102
rect 26 -106 30 -102
rect 53 -104 80 -100
rect -48 -110 37 -106
rect 53 -108 57 -104
rect 76 -108 80 -104
rect 33 -115 37 -110
rect 42 -115 46 -112
rect 61 -115 65 -112
rect -48 -119 108 -115
rect -48 -197 -44 -119
rect -38 -131 -34 -119
rect -7 -123 -3 -119
rect -23 -131 -19 -127
rect -15 -131 -11 -127
rect 1 -131 5 -127
rect -15 -135 5 -131
rect 9 -131 13 -127
rect 24 -131 28 -119
rect 42 -131 46 -119
rect 73 -123 77 -119
rect 57 -131 61 -127
rect 65 -131 69 -127
rect 81 -131 85 -127
rect 65 -135 85 -131
rect 89 -131 93 -127
rect 104 -131 108 -119
rect -41 -142 -37 -138
rect -30 -145 -26 -135
rect -7 -145 -3 -143
rect -15 -149 -3 -145
rect 16 -146 20 -135
rect 27 -143 31 -139
rect 39 -142 43 -138
rect 50 -145 54 -135
rect 73 -145 77 -143
rect -38 -165 -34 -149
rect -23 -157 -19 -153
rect -15 -157 -11 -149
rect 9 -157 13 -153
rect 1 -165 5 -161
rect 24 -165 28 -150
rect 65 -149 77 -145
rect 96 -146 100 -135
rect 111 -139 115 -94
rect 107 -143 115 -139
rect 42 -165 46 -149
rect 57 -157 61 -153
rect 65 -157 69 -149
rect 89 -157 93 -153
rect 81 -165 85 -161
rect 104 -165 108 -150
rect -38 -169 108 -165
rect -38 -173 -34 -169
rect -10 -173 -6 -169
rect 18 -173 22 -169
rect 42 -173 46 -169
rect -22 -181 -18 -177
rect 6 -181 10 -177
rect 34 -181 38 -177
rect -38 -185 -18 -181
rect -10 -185 10 -181
rect 18 -182 38 -181
rect 18 -185 43 -182
rect -38 -189 -34 -185
rect -22 -189 -18 -185
rect -10 -189 -6 -185
rect 6 -189 10 -185
rect 18 -189 22 -185
rect 34 -186 43 -185
rect 50 -184 54 -179
rect 65 -183 69 -178
rect 34 -189 38 -186
rect 76 -191 80 -177
rect -30 -197 -26 -193
rect -2 -197 2 -193
rect 26 -197 30 -193
rect 53 -195 115 -191
rect -48 -201 37 -197
rect 53 -199 57 -195
rect 76 -199 80 -195
rect 33 -207 37 -201
rect 42 -207 46 -203
rect 61 -207 65 -203
rect -48 -211 108 -207
rect -48 -289 -44 -211
rect -38 -223 -34 -211
rect -7 -215 -3 -211
rect -23 -223 -19 -219
rect -15 -223 -11 -219
rect 1 -223 5 -219
rect -15 -227 5 -223
rect 9 -223 13 -219
rect 24 -223 28 -211
rect 42 -223 46 -211
rect 73 -215 77 -211
rect 57 -223 61 -219
rect 65 -223 69 -219
rect 81 -223 85 -219
rect 65 -227 85 -223
rect 89 -223 93 -219
rect 104 -223 108 -211
rect -41 -234 -37 -230
rect -30 -237 -26 -227
rect -7 -237 -3 -235
rect -15 -241 -3 -237
rect 16 -238 20 -227
rect 27 -235 31 -231
rect 39 -234 43 -230
rect 50 -237 54 -227
rect 73 -237 77 -235
rect -38 -257 -34 -241
rect -23 -249 -19 -245
rect -15 -249 -11 -241
rect 9 -249 13 -245
rect 1 -257 5 -253
rect 24 -257 28 -242
rect 65 -241 77 -237
rect 96 -238 100 -227
rect 111 -231 115 -195
rect 107 -235 115 -231
rect 42 -257 46 -241
rect 57 -249 61 -245
rect 65 -249 69 -241
rect 89 -249 93 -245
rect 81 -257 85 -253
rect 104 -257 108 -242
rect -38 -261 108 -257
rect -38 -265 -34 -261
rect -10 -265 -6 -261
rect 18 -265 22 -261
rect 42 -265 46 -261
rect -22 -273 -18 -269
rect 6 -273 10 -269
rect 34 -273 38 -269
rect -38 -277 -18 -273
rect -10 -277 10 -273
rect 18 -274 38 -273
rect 18 -277 43 -274
rect -38 -281 -34 -277
rect -22 -281 -18 -277
rect -10 -281 -6 -277
rect 6 -281 10 -277
rect 18 -281 22 -277
rect 34 -278 43 -277
rect 50 -276 54 -271
rect 65 -275 69 -270
rect 34 -281 38 -278
rect 76 -283 80 -269
rect -30 -289 -26 -285
rect -2 -289 2 -285
rect 26 -289 30 -285
rect 53 -287 115 -283
rect -48 -293 37 -289
rect 53 -291 57 -287
rect 76 -291 80 -287
rect 33 -299 37 -293
rect 42 -299 46 -295
rect 61 -299 65 -295
rect -48 -303 108 -299
rect -48 -381 -44 -303
rect -38 -315 -34 -303
rect -7 -307 -3 -303
rect -23 -315 -19 -311
rect -15 -315 -11 -311
rect 1 -315 5 -311
rect -15 -319 5 -315
rect 9 -315 13 -311
rect 24 -315 28 -303
rect 42 -315 46 -303
rect 73 -307 77 -303
rect 57 -315 61 -311
rect 65 -315 69 -311
rect 81 -315 85 -311
rect 65 -319 85 -315
rect 89 -315 93 -311
rect 104 -315 108 -303
rect -41 -326 -37 -322
rect -30 -329 -26 -319
rect -7 -329 -3 -327
rect -15 -333 -3 -329
rect 16 -330 20 -319
rect 27 -327 31 -323
rect 39 -326 43 -322
rect 50 -329 54 -319
rect 73 -329 77 -327
rect -38 -349 -34 -333
rect -23 -341 -19 -337
rect -15 -341 -11 -333
rect 9 -341 13 -337
rect 1 -349 5 -345
rect 24 -349 28 -334
rect 65 -333 77 -329
rect 96 -330 100 -319
rect 111 -323 115 -287
rect 107 -327 115 -323
rect 42 -349 46 -333
rect 57 -341 61 -337
rect 65 -341 69 -333
rect 89 -341 93 -337
rect 81 -349 85 -345
rect 104 -349 108 -334
rect -38 -353 108 -349
rect -38 -357 -34 -353
rect -10 -357 -6 -353
rect 18 -357 22 -353
rect 42 -357 46 -353
rect -22 -365 -18 -361
rect 6 -365 10 -361
rect 34 -365 38 -361
rect -38 -369 -18 -365
rect -10 -369 10 -365
rect 18 -366 38 -365
rect 18 -369 43 -366
rect -38 -373 -34 -369
rect -22 -373 -18 -369
rect -10 -373 -6 -369
rect 6 -373 10 -369
rect 18 -373 22 -369
rect 34 -370 43 -369
rect 50 -368 54 -363
rect 65 -367 69 -362
rect 34 -373 38 -370
rect 76 -375 80 -361
rect -30 -381 -26 -377
rect -2 -381 2 -377
rect 26 -381 30 -377
rect 53 -379 80 -375
rect -48 -385 37 -381
rect 53 -383 57 -379
rect 76 -383 80 -379
rect 33 -391 37 -385
rect 42 -391 46 -387
rect 61 -391 65 -387
rect 33 -395 65 -391
<< metal2 >>
rect -23 -48 -19 -44
rect 9 -48 13 -44
rect 31 -48 35 -47
rect -23 -52 -7 -48
rect -3 -51 35 -48
rect 57 -48 61 -44
rect 89 -48 93 -44
rect -3 -52 31 -51
rect 57 -52 73 -48
rect 77 -52 93 -48
rect -19 -62 9 -58
rect 61 -62 89 -58
rect -36 -74 -30 -70
rect -36 -111 -32 -74
rect -18 -106 -14 -94
rect 10 -99 14 -94
rect 50 -99 54 -97
rect 10 -102 54 -99
rect 65 -106 69 -96
rect -18 -111 69 -106
rect -36 -114 -30 -111
rect -34 -349 -30 -114
rect -23 -139 -19 -135
rect 9 -139 13 -135
rect 31 -139 35 -138
rect -23 -143 -7 -139
rect -3 -142 35 -139
rect 57 -139 61 -135
rect 89 -139 93 -135
rect -3 -143 31 -142
rect 57 -143 73 -139
rect 77 -143 93 -139
rect -19 -153 9 -149
rect 61 -153 89 -149
rect -18 -197 -14 -185
rect 10 -190 14 -185
rect 50 -190 54 -188
rect 10 -193 54 -190
rect 65 -197 69 -187
rect -18 -202 69 -197
rect -23 -231 -19 -227
rect 9 -231 13 -227
rect 31 -231 35 -230
rect -23 -235 -7 -231
rect -3 -234 35 -231
rect 57 -231 61 -227
rect 89 -231 93 -227
rect -3 -235 31 -234
rect 57 -235 73 -231
rect 77 -235 93 -231
rect -19 -245 9 -241
rect 61 -245 89 -241
rect -18 -289 -14 -277
rect 10 -282 14 -277
rect 50 -282 54 -280
rect 10 -285 54 -282
rect 65 -289 69 -279
rect -18 -294 69 -289
rect -23 -323 -19 -319
rect 9 -323 13 -319
rect 31 -323 35 -322
rect -23 -327 -7 -323
rect -3 -326 35 -323
rect 57 -323 61 -319
rect 89 -323 93 -319
rect -3 -327 31 -326
rect 57 -327 73 -323
rect 77 -327 93 -323
rect -19 -337 9 -333
rect 61 -337 89 -333
rect -18 -381 -14 -369
rect 10 -374 14 -369
rect 50 -374 54 -372
rect 10 -377 54 -374
rect 65 -381 69 -371
rect -18 -386 69 -381
<< ntransistor >>
rect -33 -58 -31 -54
rect 21 -59 23 -55
rect 47 -58 49 -54
rect 101 -59 103 -55
rect -18 -70 -16 -66
rect -10 -70 -8 -66
rect -2 -70 0 -66
rect 6 -70 8 -66
rect 62 -70 64 -66
rect 70 -70 72 -66
rect 78 -70 80 -66
rect 86 -70 88 -66
rect -33 -86 -31 -82
rect -25 -86 -23 -82
rect -5 -86 -3 -82
rect 3 -86 5 -82
rect 23 -86 25 -82
rect 31 -86 33 -82
rect 47 -86 49 -82
rect 58 -86 60 -82
rect 73 -86 75 -82
rect -33 -149 -31 -145
rect 21 -150 23 -146
rect 47 -149 49 -145
rect 101 -150 103 -146
rect -18 -161 -16 -157
rect -10 -161 -8 -157
rect -2 -161 0 -157
rect 6 -161 8 -157
rect 62 -161 64 -157
rect 70 -161 72 -157
rect 78 -161 80 -157
rect 86 -161 88 -157
rect -33 -177 -31 -173
rect -25 -177 -23 -173
rect -5 -177 -3 -173
rect 3 -177 5 -173
rect 23 -177 25 -173
rect 31 -177 33 -173
rect 47 -177 49 -173
rect 58 -177 60 -173
rect 73 -177 75 -173
rect -33 -241 -31 -237
rect 21 -242 23 -238
rect 47 -241 49 -237
rect 101 -242 103 -238
rect -18 -253 -16 -249
rect -10 -253 -8 -249
rect -2 -253 0 -249
rect 6 -253 8 -249
rect 62 -253 64 -249
rect 70 -253 72 -249
rect 78 -253 80 -249
rect 86 -253 88 -249
rect -33 -269 -31 -265
rect -25 -269 -23 -265
rect -5 -269 -3 -265
rect 3 -269 5 -265
rect 23 -269 25 -265
rect 31 -269 33 -265
rect 47 -269 49 -265
rect 58 -269 60 -265
rect 73 -269 75 -265
rect -33 -333 -31 -329
rect 21 -334 23 -330
rect 47 -333 49 -329
rect 101 -334 103 -330
rect -18 -345 -16 -341
rect -10 -345 -8 -341
rect -2 -345 0 -341
rect 6 -345 8 -341
rect 62 -345 64 -341
rect 70 -345 72 -341
rect 78 -345 80 -341
rect 86 -345 88 -341
rect -33 -361 -31 -357
rect -25 -361 -23 -357
rect -5 -361 -3 -357
rect 3 -361 5 -357
rect 23 -361 25 -357
rect 31 -361 33 -357
rect 47 -361 49 -357
rect 58 -361 60 -357
rect 73 -361 75 -357
<< ptransistor >>
rect -18 -36 -16 -32
rect -10 -36 -8 -32
rect -2 -36 0 -32
rect 6 -36 8 -32
rect -33 -44 -31 -40
rect 62 -36 64 -32
rect 70 -36 72 -32
rect 78 -36 80 -32
rect 86 -36 88 -32
rect 21 -44 23 -40
rect 47 -44 49 -40
rect 101 -44 103 -40
rect -33 -102 -31 -98
rect -25 -102 -23 -98
rect -5 -102 -3 -98
rect 3 -102 5 -98
rect 23 -102 25 -98
rect 31 -102 33 -98
rect 47 -112 49 -108
rect 58 -112 60 -108
rect 73 -112 75 -108
rect -18 -127 -16 -123
rect -10 -127 -8 -123
rect -2 -127 0 -123
rect 6 -127 8 -123
rect -33 -135 -31 -131
rect 62 -127 64 -123
rect 70 -127 72 -123
rect 78 -127 80 -123
rect 86 -127 88 -123
rect 21 -135 23 -131
rect 47 -135 49 -131
rect 101 -135 103 -131
rect -33 -193 -31 -189
rect -25 -193 -23 -189
rect -5 -193 -3 -189
rect 3 -193 5 -189
rect 23 -193 25 -189
rect 31 -193 33 -189
rect 47 -203 49 -199
rect 58 -203 60 -199
rect 73 -203 75 -199
rect -18 -219 -16 -215
rect -10 -219 -8 -215
rect -2 -219 0 -215
rect 6 -219 8 -215
rect -33 -227 -31 -223
rect 62 -219 64 -215
rect 70 -219 72 -215
rect 78 -219 80 -215
rect 86 -219 88 -215
rect 21 -227 23 -223
rect 47 -227 49 -223
rect 101 -227 103 -223
rect -33 -285 -31 -281
rect -25 -285 -23 -281
rect -5 -285 -3 -281
rect 3 -285 5 -281
rect 23 -285 25 -281
rect 31 -285 33 -281
rect 47 -295 49 -291
rect 58 -295 60 -291
rect 73 -295 75 -291
rect -18 -311 -16 -307
rect -10 -311 -8 -307
rect -2 -311 0 -307
rect 6 -311 8 -307
rect -33 -319 -31 -315
rect 62 -311 64 -307
rect 70 -311 72 -307
rect 78 -311 80 -307
rect 86 -311 88 -307
rect 21 -319 23 -315
rect 47 -319 49 -315
rect 101 -319 103 -315
rect -33 -377 -31 -373
rect -25 -377 -23 -373
rect -5 -377 -3 -373
rect 3 -377 5 -373
rect 23 -377 25 -373
rect 31 -377 33 -373
rect 47 -387 49 -383
rect 58 -387 60 -383
rect 73 -387 75 -383
<< polycontact >>
rect -37 -51 -33 -47
rect -26 -51 -22 -47
rect 12 -52 16 -48
rect 23 -52 27 -48
rect 43 -51 47 -47
rect 54 -51 58 -47
rect 92 -52 96 -48
rect 103 -52 107 -48
rect 43 -95 47 -91
rect 54 -92 58 -88
rect 69 -91 73 -87
rect -37 -142 -33 -138
rect -26 -142 -22 -138
rect 12 -143 16 -139
rect 23 -143 27 -139
rect 43 -142 47 -138
rect 54 -142 58 -138
rect 92 -143 96 -139
rect 103 -143 107 -139
rect 43 -186 47 -182
rect 54 -183 58 -179
rect 69 -182 73 -178
rect -37 -234 -33 -230
rect -26 -234 -22 -230
rect 12 -235 16 -231
rect 23 -235 27 -231
rect 43 -234 47 -230
rect 54 -234 58 -230
rect 92 -235 96 -231
rect 103 -235 107 -231
rect 43 -278 47 -274
rect 54 -275 58 -271
rect 69 -274 73 -270
rect -37 -326 -33 -322
rect -26 -326 -22 -322
rect 12 -327 16 -323
rect 23 -327 27 -323
rect 43 -326 47 -322
rect 54 -326 58 -322
rect 92 -327 96 -323
rect 103 -327 107 -323
rect 43 -370 47 -366
rect 54 -367 58 -363
rect 69 -366 73 -362
<< ndcontact >>
rect -38 -58 -34 -54
rect -30 -58 -26 -54
rect 16 -59 20 -55
rect 24 -59 28 -55
rect 42 -58 46 -54
rect 50 -58 54 -54
rect 96 -59 100 -55
rect 104 -59 108 -55
rect -23 -70 -19 -66
rect -15 -70 -11 -66
rect 1 -70 5 -66
rect 9 -70 13 -66
rect 57 -70 61 -66
rect 65 -70 69 -66
rect 81 -70 85 -66
rect 89 -70 93 -66
rect -38 -86 -34 -82
rect -22 -86 -18 -82
rect -10 -86 -6 -82
rect 6 -86 10 -82
rect 18 -86 22 -82
rect 34 -86 38 -82
rect 42 -86 46 -82
rect 76 -86 80 -82
rect -38 -149 -34 -145
rect -30 -149 -26 -145
rect 16 -150 20 -146
rect 24 -150 28 -146
rect 42 -149 46 -145
rect 50 -149 54 -145
rect 96 -150 100 -146
rect 104 -150 108 -146
rect -23 -161 -19 -157
rect -15 -161 -11 -157
rect 1 -161 5 -157
rect 9 -161 13 -157
rect 57 -161 61 -157
rect 65 -161 69 -157
rect 81 -161 85 -157
rect 89 -161 93 -157
rect -38 -177 -34 -173
rect -22 -177 -18 -173
rect -10 -177 -6 -173
rect 6 -177 10 -173
rect 18 -177 22 -173
rect 34 -177 38 -173
rect 42 -177 46 -173
rect 76 -177 80 -173
rect -38 -241 -34 -237
rect -30 -241 -26 -237
rect 16 -242 20 -238
rect 24 -242 28 -238
rect 42 -241 46 -237
rect 50 -241 54 -237
rect 96 -242 100 -238
rect 104 -242 108 -238
rect -23 -253 -19 -249
rect -15 -253 -11 -249
rect 1 -253 5 -249
rect 9 -253 13 -249
rect 57 -253 61 -249
rect 65 -253 69 -249
rect 81 -253 85 -249
rect 89 -253 93 -249
rect -38 -269 -34 -265
rect -22 -269 -18 -265
rect -10 -269 -6 -265
rect 6 -269 10 -265
rect 18 -269 22 -265
rect 34 -269 38 -265
rect 42 -269 46 -265
rect 76 -269 80 -265
rect -38 -333 -34 -329
rect -30 -333 -26 -329
rect 16 -334 20 -330
rect 24 -334 28 -330
rect 42 -333 46 -329
rect 50 -333 54 -329
rect 96 -334 100 -330
rect 104 -334 108 -330
rect -23 -345 -19 -341
rect -15 -345 -11 -341
rect 1 -345 5 -341
rect 9 -345 13 -341
rect 57 -345 61 -341
rect 65 -345 69 -341
rect 81 -345 85 -341
rect 89 -345 93 -341
rect -38 -361 -34 -357
rect -22 -361 -18 -357
rect -10 -361 -6 -357
rect 6 -361 10 -357
rect 18 -361 22 -357
rect 34 -361 38 -357
rect 42 -361 46 -357
rect 76 -361 80 -357
<< pdcontact >>
rect -23 -36 -19 -32
rect -15 -36 -11 -32
rect -7 -36 -3 -32
rect 1 -36 5 -32
rect 9 -36 13 -32
rect -38 -44 -34 -40
rect -30 -44 -26 -40
rect 57 -36 61 -32
rect 65 -36 69 -32
rect 73 -36 77 -32
rect 81 -36 85 -32
rect 89 -36 93 -32
rect 16 -44 20 -40
rect 24 -44 28 -40
rect 42 -44 46 -40
rect 50 -44 54 -40
rect 96 -44 100 -40
rect 104 -44 108 -40
rect -38 -102 -34 -98
rect -30 -102 -26 -98
rect -22 -102 -18 -98
rect -10 -102 -6 -98
rect -2 -102 2 -98
rect 6 -102 10 -98
rect 18 -102 22 -98
rect 26 -102 30 -98
rect 34 -102 38 -98
rect 42 -112 46 -108
rect 53 -112 57 -108
rect 61 -112 65 -108
rect 76 -112 80 -108
rect -23 -127 -19 -123
rect -15 -127 -11 -123
rect -7 -127 -3 -123
rect 1 -127 5 -123
rect 9 -127 13 -123
rect -38 -135 -34 -131
rect -30 -135 -26 -131
rect 57 -127 61 -123
rect 65 -127 69 -123
rect 73 -127 77 -123
rect 81 -127 85 -123
rect 89 -127 93 -123
rect 16 -135 20 -131
rect 24 -135 28 -131
rect 42 -135 46 -131
rect 50 -135 54 -131
rect 96 -135 100 -131
rect 104 -135 108 -131
rect -38 -193 -34 -189
rect -30 -193 -26 -189
rect -22 -193 -18 -189
rect -10 -193 -6 -189
rect -2 -193 2 -189
rect 6 -193 10 -189
rect 18 -193 22 -189
rect 26 -193 30 -189
rect 34 -193 38 -189
rect 42 -203 46 -199
rect 53 -203 57 -199
rect 61 -203 65 -199
rect 76 -203 80 -199
rect -23 -219 -19 -215
rect -15 -219 -11 -215
rect -7 -219 -3 -215
rect 1 -219 5 -215
rect 9 -219 13 -215
rect -38 -227 -34 -223
rect -30 -227 -26 -223
rect 57 -219 61 -215
rect 65 -219 69 -215
rect 73 -219 77 -215
rect 81 -219 85 -215
rect 89 -219 93 -215
rect 16 -227 20 -223
rect 24 -227 28 -223
rect 42 -227 46 -223
rect 50 -227 54 -223
rect 96 -227 100 -223
rect 104 -227 108 -223
rect -38 -285 -34 -281
rect -30 -285 -26 -281
rect -22 -285 -18 -281
rect -10 -285 -6 -281
rect -2 -285 2 -281
rect 6 -285 10 -281
rect 18 -285 22 -281
rect 26 -285 30 -281
rect 34 -285 38 -281
rect 42 -295 46 -291
rect 53 -295 57 -291
rect 61 -295 65 -291
rect 76 -295 80 -291
rect -23 -311 -19 -307
rect -15 -311 -11 -307
rect -7 -311 -3 -307
rect 1 -311 5 -307
rect 9 -311 13 -307
rect -38 -319 -34 -315
rect -30 -319 -26 -315
rect 57 -311 61 -307
rect 65 -311 69 -307
rect 73 -311 77 -307
rect 81 -311 85 -307
rect 89 -311 93 -307
rect 16 -319 20 -315
rect 24 -319 28 -315
rect 42 -319 46 -315
rect 50 -319 54 -315
rect 96 -319 100 -315
rect 104 -319 108 -315
rect -38 -377 -34 -373
rect -30 -377 -26 -373
rect -22 -377 -18 -373
rect -10 -377 -6 -373
rect -2 -377 2 -373
rect 6 -377 10 -373
rect 18 -377 22 -373
rect 26 -377 30 -373
rect 34 -377 38 -373
rect 42 -387 46 -383
rect 53 -387 57 -383
rect 61 -387 65 -383
rect 76 -387 80 -383
<< m2contact >>
rect -23 -44 -19 -40
rect 9 -44 13 -40
rect 57 -44 61 -40
rect 89 -44 93 -40
rect -7 -52 -3 -48
rect 35 -51 39 -47
rect 73 -52 77 -48
rect -23 -62 -19 -58
rect 9 -62 13 -58
rect -30 -74 -26 -70
rect 57 -62 61 -58
rect 89 -62 93 -58
rect -18 -94 -14 -90
rect 10 -94 14 -90
rect 50 -97 54 -93
rect 65 -96 69 -92
rect -23 -135 -19 -131
rect 9 -135 13 -131
rect 57 -135 61 -131
rect 89 -135 93 -131
rect -7 -143 -3 -139
rect 35 -142 39 -138
rect 73 -143 77 -139
rect -23 -153 -19 -149
rect 9 -153 13 -149
rect -30 -165 -26 -161
rect 57 -153 61 -149
rect 89 -153 93 -149
rect -18 -185 -14 -181
rect 10 -185 14 -181
rect 50 -188 54 -184
rect 65 -187 69 -183
rect -23 -227 -19 -223
rect 9 -227 13 -223
rect 57 -227 61 -223
rect 89 -227 93 -223
rect -7 -235 -3 -231
rect 35 -234 39 -230
rect 73 -235 77 -231
rect -23 -245 -19 -241
rect 9 -245 13 -241
rect -30 -257 -26 -253
rect 57 -245 61 -241
rect 89 -245 93 -241
rect -18 -277 -14 -273
rect 10 -277 14 -273
rect 50 -280 54 -276
rect 65 -279 69 -275
rect -23 -319 -19 -315
rect 9 -319 13 -315
rect 57 -319 61 -315
rect 89 -319 93 -315
rect -7 -327 -3 -323
rect 35 -326 39 -322
rect 73 -327 77 -323
rect -23 -337 -19 -333
rect 9 -337 13 -333
rect -30 -349 -26 -345
rect 57 -337 61 -333
rect 89 -337 93 -333
rect -18 -369 -14 -365
rect 10 -369 14 -365
rect 50 -372 54 -368
rect 65 -371 69 -367
use 2-bitXOR 2-bitXOR_0
timestamp 1332627727
transform 1 0 14 0 1 23
box 0 0 1 1
use 2-bitXOR 2-bitXOR_1
timestamp 1332627727
transform 1 0 -27 0 1 -55
box 0 0 1 1
use 2-bitXOR 2-bitXOR_2
timestamp 1332627727
transform 1 0 53 0 1 -55
box 0 0 1 1
use 2-bitXOR 2-bitXOR_3
timestamp 1332627727
transform 1 0 -27 0 1 -146
box 0 0 1 1
use 2-bitXOR 2-bitXOR_4
timestamp 1332627727
transform 1 0 53 0 1 -146
box 0 0 1 1
use 2-bitXOR 2-bitXOR_5
timestamp 1332627727
transform 1 0 -27 0 1 -238
box 0 0 1 1
use 2-bitXOR 2-bitXOR_6
timestamp 1332627727
transform 1 0 53 0 1 -238
box 0 0 1 1
use 2-bitXOR 2-bitXOR_7
timestamp 1332627727
transform 1 0 -27 0 1 -330
box 0 0 1 1
use 2-bitXOR 2-bitXOR_8
timestamp 1332627727
transform 1 0 53 0 1 -330
box 0 0 1 1
<< labels >>
rlabel metal1 3 -76 3 -76 1 GND
rlabel metal1 -5 -27 -5 -27 5 VDD
rlabel metal1 109 -50 109 -50 7 CIN
rlabel metal1 -40 -140 -40 -140 1 A2
rlabel metal1 -39 -232 -39 -232 1 A3
rlabel metal1 -39 -325 -39 -325 1 A4
rlabel metal1 29 -141 29 -141 1 B2
rlabel metal1 29 -233 29 -233 1 B3
rlabel metal1 29 -325 29 -325 1 B4
rlabel metal1 75 -56 75 -56 1 S1
rlabel metal1 75 -147 75 -147 1 S2
rlabel metal1 75 -239 75 -239 1 S3
rlabel metal1 75 -331 75 -331 1 S4
rlabel metal1 29 -50 29 -50 1 B1
rlabel metal1 -39 -49 -39 -49 1 A1
rlabel metal1 78 -374 78 -374 1 Cout
<< end >>
