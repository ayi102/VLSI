magic
tech scmos
timestamp 1331343439
<< polysilicon >>
rect 5 24 36 26
rect 5 4 7 24
rect 18 20 20 22
rect 26 20 28 22
rect 34 20 36 24
rect 42 20 44 22
rect 5 -12 7 0
rect 5 -18 7 -16
rect 18 -27 20 16
rect 26 -27 28 16
rect 34 -27 36 16
rect 42 -27 44 16
rect 57 4 59 6
rect 57 -12 59 0
rect 18 -33 20 -31
rect 26 -35 28 -31
rect 34 -33 36 -31
rect 42 -33 44 -31
rect 57 -35 59 -16
rect 26 -37 59 -35
<< ndiffusion >>
rect 4 -16 5 -12
rect 7 -16 8 -12
rect 56 -16 57 -12
rect 59 -16 60 -12
rect 17 -31 18 -27
rect 20 -31 26 -27
rect 28 -31 29 -27
rect 33 -31 34 -27
rect 36 -31 42 -27
rect 44 -31 45 -27
<< pdiffusion >>
rect 17 16 18 20
rect 20 16 21 20
rect 25 16 26 20
rect 28 16 29 20
rect 33 16 34 20
rect 36 16 37 20
rect 41 16 42 20
rect 44 16 45 20
rect 4 0 5 4
rect 7 0 8 4
rect 56 0 57 4
rect 59 0 60 4
<< metal1 >>
rect 0 24 64 28
rect 0 4 4 24
rect 21 20 25 24
rect 13 12 17 16
rect 13 8 21 12
rect 17 4 21 8
rect 29 4 33 16
rect 37 12 41 16
rect 45 4 49 16
rect 60 4 64 24
rect 17 0 49 4
rect 8 -3 12 0
rect 52 -3 56 0
rect -3 -8 1 -4
rect 8 -7 14 -3
rect 48 -7 56 -3
rect 63 -7 67 -3
rect 8 -12 12 -7
rect 52 -12 56 -7
rect 0 -35 4 -16
rect 13 -23 49 -19
rect 13 -27 17 -23
rect 45 -27 49 -23
rect 29 -35 33 -31
rect 60 -35 64 -16
rect 0 -39 64 -35
<< metal2 >>
rect 37 -15 41 8
<< ntransistor >>
rect 5 -16 7 -12
rect 57 -16 59 -12
rect 18 -31 20 -27
rect 26 -31 28 -27
rect 34 -31 36 -27
rect 42 -31 44 -27
<< ptransistor >>
rect 18 16 20 20
rect 26 16 28 20
rect 34 16 36 20
rect 42 16 44 20
rect 5 0 7 4
rect 57 0 59 4
<< polycontact >>
rect 1 -8 5 -4
rect 14 -7 18 -3
rect 44 -7 48 -3
rect 59 -7 63 -3
<< ndcontact >>
rect 0 -16 4 -12
rect 8 -16 12 -12
rect 52 -16 56 -12
rect 60 -16 64 -12
rect 13 -31 17 -27
rect 29 -31 33 -27
rect 45 -31 49 -27
<< pdcontact >>
rect 13 16 17 20
rect 21 16 25 20
rect 29 16 33 20
rect 37 16 41 20
rect 45 16 49 20
rect 0 0 4 4
rect 8 0 12 4
rect 52 0 56 4
rect 60 0 64 4
<< m2contact >>
rect 37 8 41 12
rect 37 -19 41 -15
<< labels >>
rlabel metal1 34 -37 35 -37 1 Gnd
rlabel metal1 -2 -6 -2 -6 3 A
rlabel metal1 65 -5 65 -5 7 B
rlabel metal1 45 26 45 26 5 Vdd
rlabel metal1 40 -22 40 -22 1 Y
<< end >>
