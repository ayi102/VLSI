magic
tech scmos
timestamp 1329873755
<< polysilicon >>
rect 5 4 7 6
rect 16 4 18 6
rect 23 4 25 6
rect 39 4 41 6
rect 5 -30 7 0
rect 16 -10 18 0
rect 10 -12 18 -10
rect 10 -23 12 -12
rect 10 -25 17 -23
rect 15 -30 17 -25
rect 23 -30 25 0
rect 39 -30 41 0
rect 5 -36 7 -34
rect 15 -36 17 -34
rect 23 -36 25 -34
rect 39 -36 41 -34
<< ndiffusion >>
rect 1 -34 5 -30
rect 7 -34 10 -30
rect 14 -34 15 -30
rect 17 -34 18 -30
rect 22 -34 23 -30
rect 25 -34 26 -30
rect 38 -34 39 -30
rect 41 -34 42 -30
<< pdiffusion >>
rect 1 0 5 4
rect 7 0 16 4
rect 18 0 23 4
rect 25 0 26 4
rect 38 0 39 4
rect 41 0 42 4
<< metal1 >>
rect -3 7 43 11
rect -3 4 1 7
rect 34 4 38 7
rect -3 -7 1 -3
rect 8 -7 12 -3
rect 15 -19 19 -15
rect 26 -16 30 0
rect 26 -20 35 -16
rect 26 -23 30 -20
rect 10 -27 30 -23
rect 10 -30 14 -27
rect 26 -30 30 -27
rect 42 -30 46 0
rect -3 -37 1 -34
rect 18 -37 22 -34
rect 34 -37 38 -34
rect -3 -41 38 -37
<< ntransistor >>
rect 5 -34 7 -30
rect 15 -34 17 -30
rect 23 -34 25 -30
rect 39 -34 41 -30
<< ptransistor >>
rect 5 0 7 4
rect 16 0 18 4
rect 23 0 25 4
rect 39 0 41 4
<< polycontact >>
rect 1 -7 5 -3
rect 12 -7 16 -3
rect 19 -19 23 -15
rect 35 -20 39 -16
<< ndcontact >>
rect -3 -34 1 -30
rect 10 -34 14 -30
rect 18 -34 22 -30
rect 26 -34 30 -30
rect 34 -34 38 -30
rect 42 -34 46 -30
<< pdcontact >>
rect -3 0 1 4
rect 26 0 30 4
rect 34 0 38 4
rect 42 0 46 4
<< labels >>
rlabel metal1 2 9 2 9 4 VDD
rlabel metal1 -1 -5 -1 -5 3 A
rlabel metal1 10 -5 10 -5 1 B
rlabel metal1 2 -39 2 -39 2 GND
rlabel metal1 17 -17 17 -17 1 C
rlabel metal1 44 -18 44 -18 7 Y
<< end >>
