magic
tech scmos
timestamp 1333128998
<< polysilicon >>
rect -34 256 -9 258
rect -34 244 -32 256
rect -19 252 -17 254
rect -11 252 -9 256
rect -3 256 22 258
rect -3 252 -1 256
rect 5 252 7 254
rect -34 228 -32 240
rect -19 232 -17 248
rect -11 232 -9 248
rect -3 232 -1 248
rect 5 232 7 248
rect 20 244 22 256
rect 38 252 40 254
rect 44 252 68 254
rect 72 252 74 254
rect 38 244 40 246
rect 44 244 68 246
rect 72 244 74 246
rect -19 230 -16 232
rect -11 230 -7 232
rect -34 222 -32 224
rect -18 222 -16 230
rect -9 222 -7 230
rect -5 230 -1 232
rect 4 230 7 232
rect -5 222 -3 230
rect 4 222 6 230
rect 20 228 22 240
rect 90 236 92 238
rect 94 236 96 238
rect 111 236 113 238
rect 20 222 22 224
rect 38 221 40 223
rect 44 221 68 223
rect 72 221 74 223
rect -18 216 -16 218
rect -9 216 -7 218
rect -5 216 -3 218
rect 4 216 6 218
rect 38 213 40 215
rect 44 213 68 215
rect 72 213 74 215
rect -18 208 -16 210
rect -9 208 -7 210
rect -5 208 -3 210
rect 4 208 6 210
rect -34 202 -32 204
rect -34 186 -32 198
rect -18 196 -16 204
rect -9 196 -7 204
rect -19 194 -16 196
rect -11 194 -7 196
rect -5 196 -3 204
rect 4 196 6 204
rect 20 202 22 204
rect -5 194 -1 196
rect 4 194 7 196
rect -34 170 -32 182
rect -19 178 -17 194
rect -11 178 -9 194
rect -3 178 -1 194
rect 5 178 7 194
rect 20 186 22 198
rect 38 183 40 185
rect 44 183 68 185
rect 72 183 74 185
rect -19 172 -17 174
rect -11 170 -9 174
rect -34 168 -9 170
rect -3 170 -1 174
rect 5 172 7 174
rect 20 170 22 182
rect 90 182 92 232
rect 94 208 96 232
rect 94 206 104 208
rect 102 189 104 206
rect 111 200 113 232
rect 99 187 104 189
rect 107 198 113 200
rect 99 182 101 187
rect 107 182 109 198
rect 38 175 40 177
rect 44 175 68 177
rect 72 175 74 177
rect 90 176 92 178
rect 99 176 101 178
rect 107 176 109 178
rect -3 168 22 170
<< ndiffusion >>
rect 68 254 72 255
rect 68 246 72 252
rect -35 224 -34 228
rect -32 224 -31 228
rect 68 243 72 244
rect 89 232 90 236
rect 92 232 94 236
rect 96 232 111 236
rect 113 232 118 236
rect 19 224 20 228
rect 22 224 23 228
rect 68 223 72 224
rect -19 218 -18 222
rect -16 218 -15 222
rect -11 218 -9 222
rect -7 218 -5 222
rect -3 218 -1 222
rect 3 218 4 222
rect 6 218 7 222
rect 68 215 72 221
rect 68 212 72 213
rect -19 204 -18 208
rect -16 204 -15 208
rect -11 204 -9 208
rect -7 204 -5 208
rect -3 204 -1 208
rect 3 204 4 208
rect 6 204 7 208
rect -35 198 -34 202
rect -32 198 -31 202
rect 19 198 20 202
rect 22 198 23 202
rect 68 185 72 186
rect 68 177 72 183
rect 68 174 72 175
<< pdiffusion >>
rect -20 248 -19 252
rect -17 248 -16 252
rect -12 248 -11 252
rect -9 248 -8 252
rect -4 248 -3 252
rect -1 248 0 252
rect 4 248 5 252
rect 7 248 8 252
rect -35 240 -34 244
rect -32 240 -31 244
rect 40 254 44 255
rect 40 251 44 252
rect 40 246 44 247
rect 19 240 20 244
rect 22 240 23 244
rect 40 243 44 244
rect 40 223 44 224
rect 40 220 44 221
rect 40 215 44 216
rect 40 212 44 213
rect -35 182 -34 186
rect -32 182 -31 186
rect 19 182 20 186
rect 22 182 23 186
rect 40 185 44 186
rect 40 182 44 183
rect -20 174 -19 178
rect -17 174 -16 178
rect -12 174 -11 178
rect -9 174 -8 178
rect -4 174 -3 178
rect -1 174 0 178
rect 4 174 5 178
rect 7 174 8 178
rect 40 177 44 178
rect 89 178 90 182
rect 92 178 94 182
rect 98 178 99 182
rect 101 178 102 182
rect 106 178 107 182
rect 109 178 110 182
rect 40 174 44 175
<< metal1 >>
rect -13 262 47 266
rect -39 258 -13 259
rect -9 258 40 259
rect -39 255 40 258
rect 47 258 51 262
rect -39 244 -35 255
rect -8 252 -4 255
rect -24 244 -20 248
rect -16 245 -12 248
rect 0 245 4 248
rect -16 241 4 245
rect 8 243 12 248
rect 23 244 27 255
rect -31 236 -27 240
rect 33 243 37 255
rect 63 255 68 259
rect 63 251 67 255
rect 44 247 63 251
rect -31 232 -23 236
rect -12 233 0 237
rect 15 236 19 240
rect -31 228 -27 232
rect -8 230 -4 233
rect 11 232 19 236
rect 33 239 40 243
rect 33 235 37 239
rect -39 215 -35 224
rect -23 222 -19 225
rect -15 226 -4 230
rect -15 222 -11 226
rect 3 225 11 229
rect 7 222 11 225
rect 15 228 19 232
rect 26 231 30 235
rect 34 231 37 235
rect 33 228 37 231
rect -1 215 3 218
rect 23 215 27 224
rect -39 211 23 215
rect -39 202 -35 211
rect -15 208 -11 211
rect -31 194 -27 198
rect -23 201 -19 204
rect -23 197 -15 201
rect -1 200 3 204
rect -8 196 3 200
rect 7 201 11 204
rect 23 202 27 211
rect 33 224 40 228
rect 47 227 51 239
rect 55 235 59 240
rect 72 239 122 243
rect 33 212 37 224
rect 63 224 68 228
rect 63 220 67 224
rect 44 216 63 220
rect 33 208 40 212
rect -42 190 -38 194
rect -31 190 -23 194
rect -8 193 -4 196
rect 15 194 19 198
rect -31 186 -27 190
rect -12 189 0 193
rect 11 190 19 194
rect 26 190 29 194
rect 33 190 37 208
rect 47 194 51 209
rect 55 212 59 213
rect 75 212 79 239
rect 118 236 122 239
rect 72 208 79 212
rect 55 194 59 208
rect 75 204 79 208
rect -39 171 -35 182
rect -24 178 -20 183
rect -16 181 4 185
rect -16 178 -12 181
rect 0 178 4 181
rect 8 178 12 183
rect 15 186 19 190
rect 33 186 40 190
rect 47 189 51 190
rect -8 171 -4 174
rect 23 171 27 182
rect 33 174 37 186
rect 63 186 68 190
rect 63 182 67 186
rect 44 178 63 182
rect 33 171 40 174
rect -39 170 40 171
rect 75 174 79 200
rect 85 189 89 232
rect 103 225 107 229
rect 104 207 108 211
rect 96 196 100 203
rect 85 185 106 189
rect 85 182 89 185
rect 102 182 106 185
rect 94 174 98 178
rect 110 174 114 178
rect -39 167 37 170
rect 47 167 55 171
rect 72 170 79 174
rect 83 170 114 174
rect 33 164 37 167
rect 83 164 87 170
rect 33 160 87 164
<< metal2 >>
rect 47 243 51 262
rect 67 247 83 251
rect -24 237 -20 240
rect 8 237 12 239
rect -43 233 -16 237
rect 4 233 12 237
rect -43 206 -39 233
rect 34 231 55 235
rect -19 225 -1 229
rect 27 211 33 215
rect -46 202 -39 206
rect 29 204 33 211
rect 55 212 59 231
rect 79 229 83 247
rect 79 225 99 229
rect 107 225 111 229
rect 67 216 84 220
rect 80 212 84 216
rect 95 212 104 215
rect 80 208 99 212
rect -46 194 -42 202
rect -11 197 7 201
rect 29 200 75 204
rect 104 203 108 207
rect -24 189 -16 193
rect 4 189 12 193
rect 33 190 47 194
rect -24 187 -20 189
rect 8 187 12 189
rect 55 171 59 190
rect 80 192 96 196
rect 80 182 84 192
rect 67 178 84 182
<< ntransistor >>
rect 68 252 72 254
rect 68 244 72 246
rect -34 224 -32 228
rect 90 232 92 236
rect 94 232 96 236
rect 111 232 113 236
rect 20 224 22 228
rect -18 218 -16 222
rect -9 218 -7 222
rect -5 218 -3 222
rect 4 218 6 222
rect 68 221 72 223
rect 68 213 72 215
rect -18 204 -16 208
rect -9 204 -7 208
rect -5 204 -3 208
rect 4 204 6 208
rect -34 198 -32 202
rect 20 198 22 202
rect 68 183 72 185
rect 68 175 72 177
<< ptransistor >>
rect -19 248 -17 252
rect -11 248 -9 252
rect -3 248 -1 252
rect 5 248 7 252
rect -34 240 -32 244
rect 40 252 44 254
rect 40 244 44 246
rect 20 240 22 244
rect 40 221 44 223
rect 40 213 44 215
rect -34 182 -32 186
rect 20 182 22 186
rect 40 183 44 185
rect -19 174 -17 178
rect -11 174 -9 178
rect -3 174 -1 178
rect 5 174 7 178
rect 90 178 92 182
rect 99 178 101 182
rect 107 178 109 182
rect 40 175 44 177
<< polycontact >>
rect -13 258 -9 262
rect -23 232 -19 236
rect 47 254 51 258
rect 7 232 11 236
rect 55 240 59 244
rect 22 231 26 235
rect 47 223 51 227
rect 47 209 51 213
rect -38 190 -34 194
rect -23 190 -19 194
rect 7 190 11 194
rect 22 190 26 194
rect 47 185 51 189
rect 107 225 111 229
rect 92 199 96 203
rect 104 203 108 207
rect 47 171 51 175
<< ndcontact >>
rect 68 255 72 259
rect -39 224 -35 228
rect -31 224 -27 228
rect 68 239 72 243
rect 85 232 89 236
rect 118 232 122 236
rect 15 224 19 228
rect 23 224 27 228
rect 68 224 72 228
rect -23 218 -19 222
rect -15 218 -11 222
rect -1 218 3 222
rect 7 218 11 222
rect 68 208 72 212
rect -23 204 -19 208
rect -15 204 -11 208
rect -1 204 3 208
rect 7 204 11 208
rect -39 198 -35 202
rect -31 198 -27 202
rect 15 198 19 202
rect 23 198 27 202
rect 68 186 72 190
rect 68 170 72 174
<< pdcontact >>
rect -24 248 -20 252
rect -16 248 -12 252
rect -8 248 -4 252
rect 0 248 4 252
rect 8 248 12 252
rect -39 240 -35 244
rect -31 240 -27 244
rect 40 255 44 259
rect 40 247 44 251
rect 15 240 19 244
rect 23 240 27 244
rect 40 239 44 243
rect 40 224 44 228
rect 40 216 44 220
rect 40 208 44 212
rect -39 182 -35 186
rect -31 182 -27 186
rect 40 186 44 190
rect 15 182 19 186
rect 23 182 27 186
rect -24 174 -20 178
rect -16 174 -12 178
rect -8 174 -4 178
rect 0 174 4 178
rect 8 174 12 178
rect 40 178 44 182
rect 85 178 89 182
rect 94 178 98 182
rect 102 178 106 182
rect 110 178 114 182
rect 40 170 44 174
<< m2contact >>
rect 47 262 51 266
rect -24 240 -20 244
rect 8 239 12 243
rect 63 247 67 251
rect -16 233 -12 237
rect 0 233 4 237
rect 47 239 51 243
rect -23 225 -19 229
rect -1 225 3 229
rect 30 231 34 235
rect 23 211 27 215
rect -15 197 -11 201
rect 7 197 11 201
rect 55 231 59 235
rect 63 216 67 220
rect -46 190 -42 194
rect -16 189 -12 193
rect 0 189 4 193
rect 29 190 33 194
rect 47 190 51 194
rect 55 208 59 212
rect 55 190 59 194
rect 75 200 79 204
rect -24 183 -20 187
rect 8 183 12 187
rect 63 178 67 182
rect 99 225 103 229
rect 104 211 108 215
rect 96 192 100 196
rect 55 167 59 171
<< labels >>
rlabel metal1 -6 257 -6 257 5 VDD
rlabel metal1 -6 213 -6 213 1 GND
rlabel metal1 28 233 28 233 1 B
rlabel metal1 -11 264 -11 264 5 A
rlabel metal1 -6 191 -6 191 1 S
rlabel metal1 28 192 28 192 1 Cin
rlabel metal1 87 205 87 205 1 Cout
<< end >>
